//NOT DONE

`timescale 1ns/1ps

//transaction class
class transaction;
  
  //declare the variables for operation type
  typedef enum bit  {write = 1'b0 , read = 1'b1} oper_type;
  randc oper_type oper;
  
  //declare the other data variables
  bit rx;
  rand bit [7:0] dintx;
  bit newd;
  bit tx;
  bit [7:0] doutrx;
  bit donetx;
  bit donerx;
  
  //deep copy
  function transaction copy();
    copy = new();
    copy.rx = this.rx;
    copy.dintx = this.dintx;
    copy.newd = this.newd;
    copy.tx = this.tx;
    copy.doutrx = this.doutrx;
    copy.donetx = this.donetx;
    copy.donerx = this.donerx;
    copy.oper = this.oper;
  endfunction
  
endclass
 
//interface
interface uart_if;
  logic clk;
  logic uclktx;
  logic uclkrx;
  logic rst;
  logic rx;
  logic [7:0] dintx;
  logic newd;
  logic tx;
  logic [7:0] doutrx;
  logic donetx;
  logic donerx;
endinterface

 
//generator class
class generator;

  //declare the data variables
  transaction tr;
  mailbox #(transaction) mbx;
  event done;
  event drvnext;
  event sconext;
  int count = 0;
  
  //custom constructor
  function new(mailbox #(transaction) mbx);
    this.mbx = mbx;
    tr = new();
  endfunction
  
  //main task
  task run();
    
    repeat(count) begin
      assert(tr.randomize) else $error("[GEN] :Randomization Failed");
      mbx.put(tr.copy);
      $display("[GEN]: Oper : %0s Din : %0d",tr.oper.name(), tr.dintx);
      @(drvnext);
      @(sconext);
    end
    -> done;
    
  endtask
endclass
 
//driver class
class driver;
  
  //call the data variables
  virtual uart_if vif;
  transaction tr;
  mailbox #(transaction) mbx;
  mailbox #(bit [7:0]) mbxds;
  event drvnext;
  
  bit [7:0] din;
  bit wr = 0;  ///random operation read / write
  bit [7:0] datarx;  ///data rcvd during read
  
  //custom constructor
  function new(mailbox #(bit [7:0]) mbxds, mailbox #(transaction) mbx);
    this.mbx = mbx;
    this.mbxds = mbxds;
   endfunction
  
  //reset
  task reset();
    vif.rst <= 1'b1;
    vif.dintx <= 0;
    vif.newd <= 0;
    vif.rx <= 1'b1;
 
    repeat(5) @(posedge vif.uclktx);
    vif.rst <= 1'b0;
    @(posedge vif.uclktx);
    $display("[DRV] : RESET DONE");
    $display("----------------------------------------");
  endtask
  

  //run
  task run();
  
    forever begin
      mbx.get(tr);
      
      if(tr.oper == 1'b0)  ////data transmission
          begin
            
            @(posedge vif.uclktx);
            vif.rst <= 1'b0;
            vif.newd <= 1'b1;  ///start data sending op
            vif.rx <= 1'b1;
            vif.dintx = tr.dintx;
            @(posedge vif.uclktx);
            vif.newd <= 1'b0;
              ////wait for completion 
            //repeat(9) @(posedge vif.uclktx);
            mbxds.put(tr.dintx);
            $display("[DRV]: Data Sent : %0d", tr.dintx);
             wait(vif.donetx == 1'b1);  
             ->drvnext;  
          end
      
      else if (tr.oper == 1'b1) begin
        
                 
        @(posedge vif.uclkrx);
        vif.rst <= 1'b0;
        vif.rx <= 1'b0;
        vif.newd <= 1'b0;
        @(posedge vif.uclkrx);
                  
        for(int i=0; i<=7; i++) begin   
          @(posedge vif.uclkrx);                
          vif.rx <= $urandom;
          datarx[i] = vif.rx;                                      
        end 
                 
                 
        mbxds.put(datarx);
        
        $display("[DRV]: Data RCVD : %0d", datarx); 
        wait(vif.donerx == 1'b1);
        vif.rx <= 1'b1;
        ->drvnext;
                 
      end         
    end   
  endtask
endclass
 
 
//monitor class
class monitor;
 
  //declare the data variables
  transaction tr;
  mailbox #(bit [7:0]) mbx;
  virtual uart_if vif;

  bit [7:0] srx; //////send
  bit [7:0] rrx; ///// recv
  
  function new(mailbox #(bit [7:0]) mbx);
    this.mbx = mbx;
  endfunction
  
  task run();
    
    forever begin
      @(posedge vif.uclktx);
      if ( (vif.newd== 1'b1) && (vif.rx == 1'b1) ) begin
        
        @(posedge vif.uclktx); 
        
        ////start collecting tx data from next clock tick
        for(int i = 0; i<= 7; i++) begin 
          @(posedge vif.uclktx);
          srx[i] = vif.tx;
        end
        $display("[MON] : DATA SEND on UART TX %0d", srx);
                  
        //////////wait for done tx before proceeding next transaction        
        @(posedge vif.uclktx); 
        mbx.put(srx);
      end
      
      else if ((vif.rx == 1'b0) && (vif.newd == 1'b0) ) begin
        wait(vif.donerx == 1);
        rrx = vif.doutrx;     
        $display("[MON] : DATA RCVD RX %0d", rrx);
        @(posedge vif.uclktx); 
        mbx.put(rrx);
      end
    end  
endtask
  
 
endclass
 

//scoreboard class
class scoreboard;
  
  //declare the data variables
  mailbox #(bit [7:0]) mbxds, mbxms;
  bit [7:0] ds;
  bit [7:0] ms;
  event sconext;
  
  //custom constructor
  function new(mailbox #(bit [7:0]) mbxds, mailbox #(bit [7:0]) mbxms);
    this.mbxds = mbxds;
    this.mbxms = mbxms;
  endfunction
  
  //main task
  task run();
    forever begin
      
      mbxds.get(ds);
      mbxms.get(ms);
      
      $display("[SCO] : DRV : %0d MON : %0d", ds, ms);
      
      if(ds == ms)
        $display("DATA MATCHED");
      else
        $display("DATA MISMATCHED");
      
      $display("----------------------------------------");
      ->sconext; 
    end
  endtask
endclass
 

//environment class
class environment;
 
  generator gen;
  driver drv;
  monitor mon;
  scoreboard sco; 
  
    
  event nextgd; ///gen -> drv
  event nextgs;  /// gen -> sco
 
  mailbox #(transaction) mbxgd; ///gen - drv
  mailbox #(bit [7:0]) mbxds; /// drv - sco 
  mailbox #(bit [7:0]) mbxms;  /// mon - sco
  virtual uart_if vif;
 
  
  function new(virtual uart_if vif);
       
    mbxgd = new();
    mbxms = new();
    mbxds = new();
    
    gen = new(mbxgd);
    drv = new(mbxds,mbxgd);
    
    
 
    mon = new(mbxms);
    sco = new(mbxds, mbxms);
    
    this.vif = vif;
    drv.vif = this.vif;
    mon.vif = this.vif;
    
    gen.sconext = nextgs;
    sco.sconext = nextgs;
    
    gen.drvnext = nextgd;
    drv.drvnext = nextgd;
 
  endfunction
  
  task pre_test();
    drv.reset();
  endtask
  
  task test();
  fork
    gen.run();
    drv.run();
    mon.run();
    sco.run();
  join_any
  endtask
  
  task post_test();
    wait(gen.done.triggered);  
    $finish();
  endtask
  
  task run();
    pre_test();
    test();
    post_test();
  endtask
 
endclass
 
 
//testbench top module
module tb;
    
  uart_if vif();
  
  uarttx #(1000000, 9600) dut (vif.clk,vif.rst,vif.rx,vif.dintx,vif.newd,vif.tx,vif.doutrx,vif.donetx, vif.donerx);
  
  initial begin
    vif.clk <= 0;
  end
    
  always #10 vif.clk <= ~vif.clk;
    
  environment env;
  
  initial begin
    env = new(vif);
    env.gen.count = 5;
    env.run();
  end
      
    
  initial begin
    $dumpfile("dump.vcd");
    $dumpvars;
  end
   
  assign vif.uclktx = dut.utx.uclk;
  assign vif.uclkrx = dut.rtx.uclk;

endmodule
